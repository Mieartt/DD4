library ieee;
use ieee.std_logic_116.all
entity ammar is
port ( wednin, khcham    : in std_logic;
        fom              : out std_logic);
end entity;
architecture behavior of ammar is
